

   M<+   �������� % File created by merging: 
File1: bV 
     Linux 6.8.0-1029-azure   4 Mergecap (Wireshark) 4.4.6 (Git commit 920939a40074) 0 File created by merging: 
File1: dw 
File2: VV 
 & File created by merging: 
File1: -w 
                �      	                     �      	                     �      	                     �      	                     �      	              